package uart_pkg;

	import uvm_pkg::*;
	`include "timescale.v"	
	`include "uvm_macros.svh"
	`include "uart_xtn.sv"
	`include "uart_agt_cfg.sv"
	`include "uart_config.sv"
	`include "uart_drv.sv"
	`include "uart_monitor.sv"
	`include "uart_seqr.sv"
	`include "uart_agent.sv"
	`include "uart_seqs.sv"
	//`include "uart_v_seqr.sv"
        //`include "uart_v_seqs.sv"
	`include "uart_sb.sv"
	`include "uart_env.sv"
	`include "uart_test.sv"
endpackage 
	
